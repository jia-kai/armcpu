/*
 * $File: vga_def.vh
 * $Date: Thu Nov 28 23:25:33 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

`define VGA_ADDR_WIDTH	18
`define VGA_DATA_WIDTH	8

`define VGA_WIDTH_MULT_SHIFT 9

// vim: ft=verilog

