../simulate/02.arith_branch_prog/mem.vh