/*
 * $File: common.vh
 * $Date: Wed Nov 20 15:55:03 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

`define REGADDR_WIDTH	5
`include "cp0_def.vh"

`define SYSTEM_STARTUP_ADDR	32'h80000000

// vim: ft=verilog


