/*
 * $File: int_def.vh
 * $Date: Wed Nov 20 18:06:35 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

// definition of interrupt numbers

`define INT_TIMER	7
`define INT_PS2		6
`define INT_SERIAL	4

// vim: ft=verilog


