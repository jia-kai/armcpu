/*
 * $File: common.vh
 * $Date: Tue Nov 19 14:44:05 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

`define REGADDR_WIDTH	5
`include "cp0_regdef.vh"

// vim: ft=verilog


