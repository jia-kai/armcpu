/*
 * $File: wb_src.vh
 * $Date: Thu Nov 14 19:51:07 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

// soruce of writeback data

`define WB_SRC_WIDTH 1
`define WB_SRC_MEM	1'b0
`define WB_SRC_ALU	1'b1

// vim: ft=verilog


