/*
 * $File: multiplier_def.vh
 * $Date: Sat Nov 23 16:45:04 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

`define 

// vim: ft=verilog

