/*
 * $File: mem_opt.vh
 * $Date: Fri Nov 15 21:10:31 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */


`define MEM_OPT_WIDTH	3
`define MEM_OPT_NONE	3'b000
`define MEM_OPT_LW		3'b001
`define MEM_OPT_LBS		3'b010
`define MEM_OPT_LBU		3'b011
`define MEM_OPT_SW		3'b100
`define MEM_OPT_SB		3'b101

// vim: ft=verilog

