/*
 * $File: int_def.vh
 * $Date: Thu Nov 21 18:28:08 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

// definition of interrupt numbers

`define INT_TIMER	7
`define INT_PS2		6
`define INT_COM		4

// vim: ft=verilog


