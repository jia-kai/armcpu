../../lib/ps2_code.vh