/*
 * $File: mmu.v
 * $Date: Sat Nov 16 09:52:34 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */


// memory management unit
module mmu(
	input [31:0] read_addr);

endmodule

