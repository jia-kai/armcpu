/*
 * $File: common.vh
 * $Date: Fri Nov 15 09:55:28 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

`define REGADDR_WIDTH	5

// vim: ft=verilog


