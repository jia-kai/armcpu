../lib/flash_driver_impl.vhd