always @(*)
casex ({shift_pressed, cur_pressed})
9'bx01011010: cur_pressed_ascii = 8'hd;
9'bx00101001: cur_pressed_ascii = 8'h20;
9'bx01100110: cur_pressed_ascii = 8'h8;
9'b000011100: cur_pressed_ascii = 8'h61;
9'b100011100: cur_pressed_ascii = 8'h41;
9'b000110010: cur_pressed_ascii = 8'h62;
9'b100110010: cur_pressed_ascii = 8'h42;
9'b000100001: cur_pressed_ascii = 8'h63;
9'b100100001: cur_pressed_ascii = 8'h43;
9'b000100011: cur_pressed_ascii = 8'h64;
9'b100100011: cur_pressed_ascii = 8'h44;
9'b000100100: cur_pressed_ascii = 8'h65;
9'b100100100: cur_pressed_ascii = 8'h45;
9'b000101011: cur_pressed_ascii = 8'h66;
9'b100101011: cur_pressed_ascii = 8'h46;
9'b000110100: cur_pressed_ascii = 8'h67;
9'b100110100: cur_pressed_ascii = 8'h47;
9'b000110011: cur_pressed_ascii = 8'h68;
9'b100110011: cur_pressed_ascii = 8'h48;
9'b001000011: cur_pressed_ascii = 8'h69;
9'b101000011: cur_pressed_ascii = 8'h49;
9'b000111011: cur_pressed_ascii = 8'h6a;
9'b100111011: cur_pressed_ascii = 8'h4a;
9'b001000010: cur_pressed_ascii = 8'h6b;
9'b101000010: cur_pressed_ascii = 8'h4b;
9'b001001011: cur_pressed_ascii = 8'h6c;
9'b101001011: cur_pressed_ascii = 8'h4c;
9'b000111010: cur_pressed_ascii = 8'h6d;
9'b100111010: cur_pressed_ascii = 8'h4d;
9'b000110001: cur_pressed_ascii = 8'h6e;
9'b100110001: cur_pressed_ascii = 8'h4e;
9'b001000100: cur_pressed_ascii = 8'h6f;
9'b101000100: cur_pressed_ascii = 8'h4f;
9'b001001101: cur_pressed_ascii = 8'h70;
9'b101001101: cur_pressed_ascii = 8'h50;
9'b000010101: cur_pressed_ascii = 8'h71;
9'b100010101: cur_pressed_ascii = 8'h51;
9'b000101101: cur_pressed_ascii = 8'h72;
9'b100101101: cur_pressed_ascii = 8'h52;
9'b000011011: cur_pressed_ascii = 8'h73;
9'b100011011: cur_pressed_ascii = 8'h53;
9'b000101100: cur_pressed_ascii = 8'h74;
9'b100101100: cur_pressed_ascii = 8'h54;
9'b000111100: cur_pressed_ascii = 8'h75;
9'b100111100: cur_pressed_ascii = 8'h55;
9'b000101010: cur_pressed_ascii = 8'h76;
9'b100101010: cur_pressed_ascii = 8'h56;
9'b000011101: cur_pressed_ascii = 8'h77;
9'b100011101: cur_pressed_ascii = 8'h57;
9'b000100010: cur_pressed_ascii = 8'h78;
9'b100100010: cur_pressed_ascii = 8'h58;
9'b000110101: cur_pressed_ascii = 8'h79;
9'b100110101: cur_pressed_ascii = 8'h59;
9'b000011010: cur_pressed_ascii = 8'h7a;
9'b100011010: cur_pressed_ascii = 8'h5a;
9'b001000101: cur_pressed_ascii = 8'h30;
9'b101000101: cur_pressed_ascii = 8'h29;
9'b000010110: cur_pressed_ascii = 8'h31;
9'b100010110: cur_pressed_ascii = 8'h21;
9'b000011110: cur_pressed_ascii = 8'h32;
9'b100011110: cur_pressed_ascii = 8'h40;
9'b000100110: cur_pressed_ascii = 8'h33;
9'b100100110: cur_pressed_ascii = 8'h23;
9'b000100101: cur_pressed_ascii = 8'h34;
9'b100100101: cur_pressed_ascii = 8'h24;
9'b000101110: cur_pressed_ascii = 8'h35;
9'b100101110: cur_pressed_ascii = 8'h25;
9'b000110110: cur_pressed_ascii = 8'h36;
9'b100110110: cur_pressed_ascii = 8'h5e;
9'b000111101: cur_pressed_ascii = 8'h37;
9'b100111101: cur_pressed_ascii = 8'h26;
9'b000111110: cur_pressed_ascii = 8'h38;
9'b100111110: cur_pressed_ascii = 8'h2a;
9'b001000110: cur_pressed_ascii = 8'h39;
9'b101000110: cur_pressed_ascii = 8'h28;
default: cur_pressed_ascii = 8'b0;
endcase
