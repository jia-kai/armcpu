/*
 * $File: lohi_def.vh
 * $Date: Sat Nov 23 19:09:47 2013 +0800
 * $Author: jiakai <jia.kai66@gmail.com>
 */

`define LOHI_WRITE_OPT_WIDTH	2
`define LOHI_WRITE_NONE	2'b00
`define LOHI_WRITE_LO		2'b01
`define LOHI_WRITE_HI		2'b10

// vim: ft=verilog

